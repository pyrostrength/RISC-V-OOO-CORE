/* 
	Register status file indicating the ROB entry of 
	the instruction writing to a destination register.
	
	Indexed by respective destination register and each entry
	contains associated ROB entry.
	
	We implement register status as 2 dual port MLAB memory module 
	and 2 dual-port ALM-based memory mode
	
	For both memory modules we indicate ROB entry to which
	a destination register is assigned on next clock cycle.
	This meshes well with current system design as well as 
	accounts for corner case in which an instruction's
	source operands' register is the exact same as the 
	destination register.
	
	regCommit is destination register of currently committing instruction.
	regCommit is only relevant for busy buffers.
	destROB is ROB entry writing to a destination register.
	destReg is destination register.
	
	Write enable is active if instruction writes to a
	destination register. If destination register
	is x0 value to be passed is changed to zero.
	
	destRegD is destReg in decode stage,destRegF is destReg in
	write RS stage.
	
*/


module register_status #(parameter REG = 4, DEPTH = 31, ROB = 2, WIDTH = 31)
								(input logic clk,we,
								 input logic[REG:0] rs1,rs2,destRegD,regCommit,destRegW,
								 input logic[ROB:0] destROB, // ROB entry that writes to a destination register.
								 output logic[ROB:0] rob1,rob2,
								 output logic[WIDTH:0] regStatusSnap,
								 output logic busy1,busy2); //rob1 and rob2 are {valid,ROB entry}
							 
							 
							   /*Two dual port MLAB memory modules
								storing ROB entry associated with
								specific register */
								
								logic[ROB:0] src1ROB[0:DEPTH];
								
								logic[ROB:0] src2ROB[0:DEPTH];
								
								logic[WIDTH:0] busyVectorI,busyVectorF;
								
								/*
								For instruction in decode stage,we 
								occupy it's destination register in the rename
								stage where we have ROB entry the instruction
								occupies*/
								
								/*Write control logic that sorts out
								destination register of current instruction
								and register of committing instruction.
								Indicate busyness of register in decode
								stage but mark ROB entry associated with
								instruction in rename stage*/
								always_comb begin
									busyVectorI = busyVectorF;
									if(destRegD != regCommit) begin
										busyVectorI[destRegD] = 1'b1;
										busyVectorI[regCommit] = 1'b0;
									end
									if(destRegD == regCommit) begin
										busyVectorI[destRegD] = 1'b1;
									end
								end
								
								/*Sorts out producing the relevant busy signals for
								instruction source operands and register status
								snapshot*/
								always_comb begin
									busy1 = (regCommit == rs1)  ? 1'b0 : busyVectorF[rs1];
									busy2 = (regCommit == rs2) ? 1'b0 : busyVectorF[rs2];
									regStatusSnap = busyVectorF;
								end
									
								/*Provide for asynchrnous read with new data
								behaviour on read during write to account for
								case in which an instruction in rename stage indicates
								its dependency*/
								always_comb begin
									rob1 = src1ROB[rs1];
									rob2 = src2ROB[rs2];
								end
									
								/* Sequential write on positive clock edge*/
								always @(posedge clk) begin
									if(we) begin
											src1ROB[destRegW] <= destROB;
											src2ROB[destRegW] <= destROB;
									end
									busyVectorF <= busyVectorI;
								end			
																
endmodule